module A;

logic a;

always_comb begin
    a = b | c;
end

endmodule
